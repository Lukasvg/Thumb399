
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

package MemoryInit is
  type mem is array(0 to 150) of std_logic_vector(7 downto 0);
  type register_file_t is array(0 to 15) of unsigned(31 downto 0);
  function InitializeMemory return mem;
  function RamSetup return register_file_t;
end;

package body MemoryInit is 
  -- Registers R0-R15 Registers Cleared
  function RamSetup return register_file_t is 
    variable temp : register_file_t;
  begin
    temp(0) := "00000000000000000000000000000000";
    temp(1) := "00000000000000000000000000000000";
    temp(2) := "00000000000000000000000000000000"; 
    temp(3) := "00000000000000000000000000000000";
    temp(4) := "00000000000000000000000000000000";
    temp(5) := "00000000000000000000000000000000";
    temp(6) := "00000000000000000000000000000000";
    temp(7) := "00000000000000000000000000000000";
    temp(8) := "00000000000000000000000000000000";
    temp(9) := "00000000000000000000000000000000";
    temp(10):= "00000000000000000000000000000000";
    temp(11):= "00000000000000000000000000000000";
    temp(12):= "00000000000000000000000000000000";
    temp(13):= "00000000000000000000000000000000";
    temp(14):= "00000000000000000000000000000000";
    temp(15):= "00000000000000000000000000000000";
    return temp;
  end function; 	 
 	 
 	-- Memory initialization function required
  function InitializeMemory return mem is
    variable temp: mem;
  begin
    -- MOV R0, #2 -------------
    -- 1st Half 1st Instruction
    temp(0) := "00100" & "000";
    -- 2nd Half 1st Instruction
    temp(1) := "00000010";
    ----------------------------
    -- MOV R1, R0 --------------
    temp(2) := "01000110";
    temp(3) := "0" & "0000" & "001";
    ---------------------------
    -- MOV R9, R1 --------------
    temp(4) := "01000110";
    temp(5) := "1" & "0001" & "001";  
    ----------------------------
    -- ASR R2, R1, #4 ----------
    temp(6) := "00010" & "001";
    temp(7) := "00" & "001" & "010"; 
    ----------------------------
    -- MOV R1, #2 --------------
    temp(8) := "00100" & "001";
    temp(9) := "00000010"; 
    ----------------------------
    -- MOV R2, #4 --------------
    temp(10) := "00100" & "010";
    temp(11) := "00000100"; 
    ----------------------------
    -- ASR R2, R1 --------------
    temp(12) := "01000001";
    temp(13) := "00" & "001" & "010"; 
    ----------------------------
    -- ADD R1, #11 -------------
    temp(14) := "00110" & "001";
    temp(15) := "00001011"; 
    ----------------------------
    -- Add R3, R2, R1 -- Add Registers
    temp(16) := "0001100" & "0";
    temp(17) := "01" & "010" & "011";  
    ----------------------------
    -- ADD R8, R4 --------------
    temp(18) := "01000100"; 
    temp(19) := "1" & "0001" & "000"; 
    ----------------------------
    
    -- Add Stack Pointer
    -- Clear Stack Pointer
    -- MOV R1, #0 --------------
    temp(20) := "00100" & "001";
    temp(21) := "00000000";
    ----------------------------
    -- MOV R13, R1 -------------
    temp(22) := "01000110"; 
    temp(23) := "1" & "0001" & "101";  
    ----------------------------
    -- Add R1, #2 --------------
    temp(24) := "10101" & "001";
    temp(25) := "00000010"; 
    ----------------------------
    -- Add #1 , SP -------------
    temp(26) := "10110000";
    temp(27) := "0" & "0000001"; 
    ----------------------------

    -- PC Addition
    -- MOV R1, #0 --------------
    temp(28) := "00100" & "001";
    temp(29) := "00000000"; 
    ----------------------------
    -- ADD R1, #1 --------------
    temp(30) := "10100" & "001";
    temp(31) := "00000001"; 
    ----------------------------

    -- ADD With Carry
    -- MOV R1, #32 -------------
    temp(32) := "00100" & "001";
    temp(33) := "00011111"; 
    ----------------------------
    -- MOV R2, #1 --------------
    temp(34) := "00100" & "010";
    temp(35) := "00000001"; 
    ----------------------------
    -- MOV R3, #1 --------------
    temp(36) := "00100" & "011";
    temp(37) := "00000001"; 
    ----------------------------
    -- LSL R2, R1 --------------
    temp(38) := "01000000";
    temp(39) := "10" & "001" & "010"; 
    ----------------------------
    -- LSL R3, R1 --------------
    temp(40) := "01000000";
    temp(41) := "10" & "001" & "011"; 
    ----------------------------
     -- Add R3, R2, R3 ---------
    temp(42) := "0001100" & "0";
    temp(43) := "11" & "010" & "011";
    ----------------------------
    -- ADC R3, R2 -- With Carry-
    temp(44) := "01000001";
    temp(45) := "01" & "010" & "011";     
    ----------------------------
    
    --LSL Instructions
    -- MOV R1, #1 --------------
    temp(46) := "00100" & "001";
    temp(47) := "00000001"; 
    ----------------------------
    -- LSL R2, R1, #4 ----------
    temp(48) := "00000" & "001";
    temp(49) := "00" & "001" & "010"; 
    ----------------------------
    
    --LSL Register
    -- MOV R1, #4 --------------
    temp(50) := "00100" & "001";
    temp(51) := "00000100"; 
    ----------------------------
    -- MOV R2, #1 --------------
    temp(52) := "00100" & "010";
    temp(53) := "00000001"; 
    ----------------------------
    
    -- LSL R2, R1 --------------
    temp(54) := "01000000";
    temp(55) := "10" & "001" & "010"; 
    ----------------------------
    -- LSR R2, R1, #4 ----------
    temp(56) := "00001" & "001";
    temp(57) := "00" & "001" & "010"; 
    ----------------------------
    
    -- MOV R1, #4---------------
    temp(58) := "00100" & "001"; 
    temp(59) := "00000100";
    ----------------------------
    -- MOV R2, #16--------------
    temp(60) := "00100" & "010"; 
    temp(61) := "00010000";
    ----------------------------
    -- LSR R2, R1 --------------
    temp(62) := "01000000";
    temp(63) := "11" & "001" & "010"; 
    ----------------------------
    
    -- ROR
    -- MOV R1, #4 --------------
    temp(64) := "00100" & "001"; 
    temp(65) := "00000100"; 
    ----------------------------
    -- MOV R2, #16 -------------
    temp(66) := "00100" & "010";
 
  temp(67) := "00010000"; 
    ----------------------------
    -- ROR R2, R1---------------
    temp(68) := "01000001";
   
temp(69) :="11" & "001" & "010"; 
    ----------------------------
    
    -- Immediate Add
    -- MOV R0, #0 --------------
    temp(70) := "00100" & "000"; 
    temp(71) := "00000000"; 
    ----------------------------
    -- MOV R1, #0 --------------
    temp(72) := "00100" & "001";
    temp(73) := "00000000"; 
    ----------------------------
    -- ADD R1, R0, #1 ----------
    temp(74) := "0001110" & "0";
    temp(75) := "01" & "000" & "001"; 
    ----------------------------
    -- ADD R2, R1, #5 ----------
    temp(76) := "0001110" & "1";
    temp(77) := "01" & "001" & "010";
    ----------------------------
    -- ADD R3, R2, #7 ----------
    temp(78) := "0001110" & "1";
    temp(79) := "11" & "010" & "011"; 
    ----------------------------
    
    -- ADD IMM8
    -- MOV R1, #0 --------------
    temp(80) := "00100" & "001";
    temp(81) := "00000000";
    ---------------------------- 
    -- MOV R8, R1 --------------
    temp(82) := "01000110"; 
    temp(83) := "1" & "0001" & "000"; 
    ----------------------------
    -- MOV R4, #1 --------------
    temp(84) := "00100" & "100";
    temp(85) := "00000001"; 
    ----------------------------
    -- ADD R1, #11 -------------
    temp(86) := "00110" & "001";
   
 temp(87) := "00001011"; 
   
 ---------------------------
   
 
  
 -- Logical Operations
  
 -- MOV R1, #32 -------------
    temp(88) := "00100" & "001";
    temp(89) := "00011111"; 
    ----------------------------
    -- MOV R2, #32 -------------
    temp(90) := "00100" & "010";
    temp(91) := "00011111"; 
    ----------------------------
    -- AND R2, R1 --------------
    temp(92) := "01000000";
    temp(93) := "00" & "001" & "010"; 
    ----------------------------
    -- BIC R2, R1 --------------
    temp(94) := "01000011";
    temp(95) := "10" & "001" & "010"; 
    ----------------------------
    -- EOR R2, R1 --------------
    temp(96) := "01000000";
    temp(97) := "01" & "001" & "010"; 
    ----------------------------
    -- MVN R2, R1 --------------
    temp(98) := "01000011";
    temp(99) := "11" & "001" & "010";
    ---------------------------- 
    -- MOV R1, #32 -------------
    temp(100) := "00100" & "001";
    temp(101) := "00011111"; 
    ----------------------------
    -- MOV R2, #63 -------------
    temp(102) := "00100" & "010"; 
    temp(103) := "00111111";
    ----------------------------
    -- OR R2, R1 ---------------
    temp(104) := "01000011";
    temp(105) := "00" & "001" & "010"; 
    ----------------------------
    
    -- Branching Operations
    -- MOV R1, #4 --------------
    temp(106) := "00100" & "001";
    temp(107) := "00000100";
    ----------------------------
    -- B + 4 -------------------
    temp(108) := "11100" & "000";
    temp(109) := "00000110";
    ----------------------------
    --ADD R1, #2 ---------------
    temp(114) := "00110" & "001";
    temp(115) := "00000010";
    ----------------------------
    
    -- MOV R0, #4 --------------
    temp(116) := "00100" & "000";
    temp(117) := "01111010";
    ----------------------------
    -- BX R0 -------------------
    temp(118) := "010001" & "11";
    temp(119) := "0" & "0000" & "000";
    ----------------------------
    --ADD R1, #2 ---------------
    temp(122) := "00110" & "001";
    temp(123) := "00000010";
    ----------------------------
    
    -- MOV R0, #4 --------------
    temp(124) := "00100" & "000";
    temp(125) := "10000010";
    ----------------------------
    -- BLX R0 ------------------
    temp(126) := "010001" & "11";
    temp(127) := "1" & "0000" & "000";
    ----------------------------
    --ADD R1, #2 ---------------
    temp(130) := "00110" & "001";
    temp(131) := "00000010";
    ----------------------------
    
    -- BL + 10 -----------------
    temp(132) := "11110" & "0" & "00";
    temp(133) := "00000000";
    temp(134) := "11" & "1" & "1" & "1" & "000";
    temp(135) := "01000110";
    ---------------------------
    --ADD R1, #2 ---------------
    temp(140) := "00110" & "001";
    temp(141) := "00000010";
    ----------------------------
    
    
    return temp;
  end function;
end package body;